module memCtrl(
    input clk,
    input rst,
    input rdy
);

endmodule