module register(
    input clk,
    input rst,
    input rdy
);

endmodule